** Profile: "System_Decoder-first"  [ D:\Orcad\lab1\first-pspicefiles\system_decoder\first.sim ] 

** Creating circuit file "first.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.INC "../../../text1.inc" 
.STMLIB "D:/Orcad/signals/reset.stl" 
.STMLIB "../../../first-pspicefiles/first.stl" 
* From [PSPICE NETLIST] section of C:\Users\bohda\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN/OP  0 10us 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\System_Decoder.net" 


.END
