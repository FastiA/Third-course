** Profile: "SCHEMATIC1-MonteCarlo"  [ D:\Orcad\lab4\amplif-pspicefiles\schematic1\montecarlo.sim ] 

** Creating circuit file "MonteCarlo.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../amplif-pspicefiles/amplif.lib" 
* From [PSPICE NETLIST] section of C:\Users\bohda\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC LIN 20 90k 110k
.WCASE AC V([[Out]]) YMAX RANGE(90k,110k)  OUTPUT ALL VARY DEV  HI 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
