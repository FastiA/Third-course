** Profile: "SCHEMATIC1-ACsweep"  [ D:\Orcad\lab2\lab2-pspicefiles\schematic1\acsweep.sim ] 

** Creating circuit file "ACsweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "D:\Orcad\lab2\lab2-pspicefiles\schematic1\ACsweep\ACsweep_profile.inc" 
* Local Libraries :
.INC "../../../clip.inc" 
* From [PSPICE NETLIST] section of C:\Users\bohda\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 11 10 100Meg
.NOISE V([OUT]) V_Vin 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
