** Profile: "SCHEMATIC1-WorstCase"  [ D:\Orcad\lab4\chebishev-pspicefiles\schematic1\worstcase.sim ] 

** Creating circuit file "WorstCase.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../chebishev-pspicefiles/chebishev.lib" 
* From [PSPICE NETLIST] section of C:\Users\bohda\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 50 100 1Meg
.WCASE AC V([OUT]) YMAX  OUTPUT ALL VARY DEV  HI DEVICES RC 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
