** Profile: "SCHEMATIC1-dcsweep"  [ D:\Orcad\lab2\lab2-pspicefiles\schematic1\dcsweep.sim ] 

** Creating circuit file "dcsweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "D:\Orcad\lab2\lab2-pspicefiles\schematic1\dcsweep\dcsweep_profile.inc" 
* Local Libraries :
.INC "../../../clip.inc" 
* From [PSPICE NETLIST] section of C:\Users\bohda\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC TEMP LIST 0 25 75 125  
+ LIN V_Vin -5 5 1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
